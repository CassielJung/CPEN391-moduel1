// step4.v

// Generated using ACDS version 19.1 670

`timescale 1 ps / 1 ps
module step4 (
		input  wire       clk_clk,       //   clk.clk
		output wire [6:0] hex0_export,   //  hex0.export
		output wire [6:0] hex1_export,   //  hex1.export
		output wire [6:0] hex2_export,   //  hex2.export
		output wire [6:0] hex3_export,   //  hex3.export
		output wire [6:0] hex4_export,   //  hex4.export
		output wire [6:0] hex5_export,   //  hex5.export
		output wire [9:0] ledr_export,   //  ledr.export
		input  wire       reset_reset_n, // reset.reset_n
		input  wire [9:0] sw_export      //    sw.export
	);

	wire  [31:0] nios2_processor_data_master_readdata;                          // mm_interconnect_0:nios2_processor_data_master_readdata -> nios2_processor:d_readdata
	wire         nios2_processor_data_master_waitrequest;                       // mm_interconnect_0:nios2_processor_data_master_waitrequest -> nios2_processor:d_waitrequest
	wire         nios2_processor_data_master_debugaccess;                       // nios2_processor:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_processor_data_master_debugaccess
	wire  [18:0] nios2_processor_data_master_address;                           // nios2_processor:d_address -> mm_interconnect_0:nios2_processor_data_master_address
	wire   [3:0] nios2_processor_data_master_byteenable;                        // nios2_processor:d_byteenable -> mm_interconnect_0:nios2_processor_data_master_byteenable
	wire         nios2_processor_data_master_read;                              // nios2_processor:d_read -> mm_interconnect_0:nios2_processor_data_master_read
	wire         nios2_processor_data_master_readdatavalid;                     // mm_interconnect_0:nios2_processor_data_master_readdatavalid -> nios2_processor:d_readdatavalid
	wire         nios2_processor_data_master_write;                             // nios2_processor:d_write -> mm_interconnect_0:nios2_processor_data_master_write
	wire  [31:0] nios2_processor_data_master_writedata;                         // nios2_processor:d_writedata -> mm_interconnect_0:nios2_processor_data_master_writedata
	wire  [31:0] nios2_processor_instruction_master_readdata;                   // mm_interconnect_0:nios2_processor_instruction_master_readdata -> nios2_processor:i_readdata
	wire         nios2_processor_instruction_master_waitrequest;                // mm_interconnect_0:nios2_processor_instruction_master_waitrequest -> nios2_processor:i_waitrequest
	wire  [18:0] nios2_processor_instruction_master_address;                    // nios2_processor:i_address -> mm_interconnect_0:nios2_processor_instruction_master_address
	wire         nios2_processor_instruction_master_read;                       // nios2_processor:i_read -> mm_interconnect_0:nios2_processor_instruction_master_read
	wire         nios2_processor_instruction_master_readdatavalid;              // mm_interconnect_0:nios2_processor_instruction_master_readdatavalid -> nios2_processor:i_readdatavalid
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;      // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;        // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest;     // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;         // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;            // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;           // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;       // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire  [31:0] mm_interconnect_0_nios2_processor_debug_mem_slave_readdata;    // nios2_processor:debug_mem_slave_readdata -> mm_interconnect_0:nios2_processor_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_processor_debug_mem_slave_waitrequest; // nios2_processor:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_processor_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_processor_debug_mem_slave_debugaccess; // mm_interconnect_0:nios2_processor_debug_mem_slave_debugaccess -> nios2_processor:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_processor_debug_mem_slave_address;     // mm_interconnect_0:nios2_processor_debug_mem_slave_address -> nios2_processor:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_processor_debug_mem_slave_read;        // mm_interconnect_0:nios2_processor_debug_mem_slave_read -> nios2_processor:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_processor_debug_mem_slave_byteenable;  // mm_interconnect_0:nios2_processor_debug_mem_slave_byteenable -> nios2_processor:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_processor_debug_mem_slave_write;       // mm_interconnect_0:nios2_processor_debug_mem_slave_write -> nios2_processor:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_processor_debug_mem_slave_writedata;   // mm_interconnect_0:nios2_processor_debug_mem_slave_writedata -> nios2_processor:debug_mem_slave_writedata
	wire         mm_interconnect_0_onchip_memory_s1_chipselect;                 // mm_interconnect_0:onchip_memory_s1_chipselect -> onchip_memory:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory_s1_readdata;                   // onchip_memory:readdata -> mm_interconnect_0:onchip_memory_s1_readdata
	wire  [14:0] mm_interconnect_0_onchip_memory_s1_address;                    // mm_interconnect_0:onchip_memory_s1_address -> onchip_memory:address
	wire   [3:0] mm_interconnect_0_onchip_memory_s1_byteenable;                 // mm_interconnect_0:onchip_memory_s1_byteenable -> onchip_memory:byteenable
	wire         mm_interconnect_0_onchip_memory_s1_write;                      // mm_interconnect_0:onchip_memory_s1_write -> onchip_memory:write
	wire  [31:0] mm_interconnect_0_onchip_memory_s1_writedata;                  // mm_interconnect_0:onchip_memory_s1_writedata -> onchip_memory:writedata
	wire         mm_interconnect_0_onchip_memory_s1_clken;                      // mm_interconnect_0:onchip_memory_s1_clken -> onchip_memory:clken
	wire         mm_interconnect_0_timer_s1_chipselect;                         // mm_interconnect_0:timer_s1_chipselect -> timer:chipselect
	wire  [15:0] mm_interconnect_0_timer_s1_readdata;                           // timer:readdata -> mm_interconnect_0:timer_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_s1_address;                            // mm_interconnect_0:timer_s1_address -> timer:address
	wire         mm_interconnect_0_timer_s1_write;                              // mm_interconnect_0:timer_s1_write -> timer:write_n
	wire  [15:0] mm_interconnect_0_timer_s1_writedata;                          // mm_interconnect_0:timer_s1_writedata -> timer:writedata
	wire         mm_interconnect_0_hex5_s1_chipselect;                          // mm_interconnect_0:HEX5_s1_chipselect -> HEX5:chipselect
	wire  [31:0] mm_interconnect_0_hex5_s1_readdata;                            // HEX5:readdata -> mm_interconnect_0:HEX5_s1_readdata
	wire   [1:0] mm_interconnect_0_hex5_s1_address;                             // mm_interconnect_0:HEX5_s1_address -> HEX5:address
	wire         mm_interconnect_0_hex5_s1_write;                               // mm_interconnect_0:HEX5_s1_write -> HEX5:write_n
	wire  [31:0] mm_interconnect_0_hex5_s1_writedata;                           // mm_interconnect_0:HEX5_s1_writedata -> HEX5:writedata
	wire         mm_interconnect_0_hex4_s1_chipselect;                          // mm_interconnect_0:HEX4_s1_chipselect -> HEX4:chipselect
	wire  [31:0] mm_interconnect_0_hex4_s1_readdata;                            // HEX4:readdata -> mm_interconnect_0:HEX4_s1_readdata
	wire   [1:0] mm_interconnect_0_hex4_s1_address;                             // mm_interconnect_0:HEX4_s1_address -> HEX4:address
	wire         mm_interconnect_0_hex4_s1_write;                               // mm_interconnect_0:HEX4_s1_write -> HEX4:write_n
	wire  [31:0] mm_interconnect_0_hex4_s1_writedata;                           // mm_interconnect_0:HEX4_s1_writedata -> HEX4:writedata
	wire         mm_interconnect_0_hex3_s1_chipselect;                          // mm_interconnect_0:HEX3_s1_chipselect -> HEX3:chipselect
	wire  [31:0] mm_interconnect_0_hex3_s1_readdata;                            // HEX3:readdata -> mm_interconnect_0:HEX3_s1_readdata
	wire   [1:0] mm_interconnect_0_hex3_s1_address;                             // mm_interconnect_0:HEX3_s1_address -> HEX3:address
	wire         mm_interconnect_0_hex3_s1_write;                               // mm_interconnect_0:HEX3_s1_write -> HEX3:write_n
	wire  [31:0] mm_interconnect_0_hex3_s1_writedata;                           // mm_interconnect_0:HEX3_s1_writedata -> HEX3:writedata
	wire         mm_interconnect_0_hex2_s1_chipselect;                          // mm_interconnect_0:HEX2_s1_chipselect -> HEX2:chipselect
	wire  [31:0] mm_interconnect_0_hex2_s1_readdata;                            // HEX2:readdata -> mm_interconnect_0:HEX2_s1_readdata
	wire   [1:0] mm_interconnect_0_hex2_s1_address;                             // mm_interconnect_0:HEX2_s1_address -> HEX2:address
	wire         mm_interconnect_0_hex2_s1_write;                               // mm_interconnect_0:HEX2_s1_write -> HEX2:write_n
	wire  [31:0] mm_interconnect_0_hex2_s1_writedata;                           // mm_interconnect_0:HEX2_s1_writedata -> HEX2:writedata
	wire         mm_interconnect_0_hex1_s1_chipselect;                          // mm_interconnect_0:HEX1_s1_chipselect -> HEX1:chipselect
	wire  [31:0] mm_interconnect_0_hex1_s1_readdata;                            // HEX1:readdata -> mm_interconnect_0:HEX1_s1_readdata
	wire   [1:0] mm_interconnect_0_hex1_s1_address;                             // mm_interconnect_0:HEX1_s1_address -> HEX1:address
	wire         mm_interconnect_0_hex1_s1_write;                               // mm_interconnect_0:HEX1_s1_write -> HEX1:write_n
	wire  [31:0] mm_interconnect_0_hex1_s1_writedata;                           // mm_interconnect_0:HEX1_s1_writedata -> HEX1:writedata
	wire         mm_interconnect_0_hex0_s1_chipselect;                          // mm_interconnect_0:HEX0_s1_chipselect -> HEX0:chipselect
	wire  [31:0] mm_interconnect_0_hex0_s1_readdata;                            // HEX0:readdata -> mm_interconnect_0:HEX0_s1_readdata
	wire   [1:0] mm_interconnect_0_hex0_s1_address;                             // mm_interconnect_0:HEX0_s1_address -> HEX0:address
	wire         mm_interconnect_0_hex0_s1_write;                               // mm_interconnect_0:HEX0_s1_write -> HEX0:write_n
	wire  [31:0] mm_interconnect_0_hex0_s1_writedata;                           // mm_interconnect_0:HEX0_s1_writedata -> HEX0:writedata
	wire         mm_interconnect_0_ledr_s1_chipselect;                          // mm_interconnect_0:LEDR_s1_chipselect -> LEDR:chipselect
	wire  [31:0] mm_interconnect_0_ledr_s1_readdata;                            // LEDR:readdata -> mm_interconnect_0:LEDR_s1_readdata
	wire   [1:0] mm_interconnect_0_ledr_s1_address;                             // mm_interconnect_0:LEDR_s1_address -> LEDR:address
	wire         mm_interconnect_0_ledr_s1_write;                               // mm_interconnect_0:LEDR_s1_write -> LEDR:write_n
	wire  [31:0] mm_interconnect_0_ledr_s1_writedata;                           // mm_interconnect_0:LEDR_s1_writedata -> LEDR:writedata
	wire  [31:0] mm_interconnect_0_sw_s1_readdata;                              // SW:readdata -> mm_interconnect_0:SW_s1_readdata
	wire   [1:0] mm_interconnect_0_sw_s1_address;                               // mm_interconnect_0:SW_s1_address -> SW:address
	wire         irq_mapper_receiver0_irq;                                      // jtag_uart:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                      // timer:irq -> irq_mapper:receiver1_irq
	wire  [31:0] nios2_processor_irq_irq;                                       // irq_mapper:sender_irq -> nios2_processor:irq
	wire         rst_controller_reset_out_reset;                                // rst_controller:reset_out -> [HEX0:reset_n, HEX1:reset_n, HEX2:reset_n, HEX3:reset_n, HEX4:reset_n, HEX5:reset_n, LEDR:reset_n, SW:reset_n, jtag_uart:rst_n, mm_interconnect_0:jtag_uart_reset_reset_bridge_in_reset_reset]
	wire         rst_controller_001_reset_out_reset;                            // rst_controller_001:reset_out -> [irq_mapper:reset, mm_interconnect_0:nios2_processor_reset_reset_bridge_in_reset_reset, nios2_processor:reset_n, onchip_memory:reset, rst_translator:in_reset, timer:reset_n]
	wire         rst_controller_001_reset_out_reset_req;                        // rst_controller_001:reset_req -> [nios2_processor:reset_req, onchip_memory:reset_req, rst_translator:reset_req_in]
	wire         nios2_processor_debug_reset_request_reset;                     // nios2_processor:debug_reset_request -> rst_controller_001:reset_in1

	step4_HEX0 hex0 (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_hex0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex0_s1_readdata),   //                    .readdata
		.out_port   (hex0_export)                           // external_connection.export
	);

	step4_HEX0 hex1 (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_hex1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex1_s1_readdata),   //                    .readdata
		.out_port   (hex1_export)                           // external_connection.export
	);

	step4_HEX0 hex2 (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_hex2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex2_s1_readdata),   //                    .readdata
		.out_port   (hex2_export)                           // external_connection.export
	);

	step4_HEX0 hex3 (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_hex3_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex3_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex3_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex3_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex3_s1_readdata),   //                    .readdata
		.out_port   (hex3_export)                           // external_connection.export
	);

	step4_HEX0 hex4 (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_hex4_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex4_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex4_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex4_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex4_s1_readdata),   //                    .readdata
		.out_port   (hex4_export)                           // external_connection.export
	);

	step4_HEX0 hex5 (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_hex5_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex5_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex5_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex5_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex5_s1_readdata),   //                    .readdata
		.out_port   (hex5_export)                           // external_connection.export
	);

	step4_LEDR ledr (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_ledr_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_ledr_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_ledr_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_ledr_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_ledr_s1_readdata),   //                    .readdata
		.out_port   (ledr_export)                           // external_connection.export
	);

	step4_SW sw (
		.clk      (clk_clk),                          //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),  //               reset.reset_n
		.address  (mm_interconnect_0_sw_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_sw_s1_readdata), //                    .readdata
		.in_port  (sw_export)                         // external_connection.export
	);

	step4_jtag_uart jtag_uart (
		.clk            (clk_clk),                                                   //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                   //               irq.irq
	);

	step4_nios2_processor nios2_processor (
		.clk                                 (clk_clk),                                                       //                       clk.clk
		.reset_n                             (~rst_controller_001_reset_out_reset),                           //                     reset.reset_n
		.reset_req                           (rst_controller_001_reset_out_reset_req),                        //                          .reset_req
		.d_address                           (nios2_processor_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_processor_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_processor_data_master_read),                              //                          .read
		.d_readdata                          (nios2_processor_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_processor_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_processor_data_master_write),                             //                          .write
		.d_writedata                         (nios2_processor_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                     (nios2_processor_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (nios2_processor_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_processor_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_processor_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_processor_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_processor_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (nios2_processor_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (nios2_processor_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_processor_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_processor_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_processor_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_processor_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_processor_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_processor_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_processor_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_processor_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_processor_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                               // custom_instruction_master.readra
	);

	step4_onchip_memory onchip_memory (
		.clk        (clk_clk),                                       //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory_s1_byteenable), //       .byteenable
		.reset      (rst_controller_001_reset_out_reset),            // reset1.reset
		.reset_req  (rst_controller_001_reset_out_reset_req),        //       .reset_req
		.freeze     (1'b0)                                           // (terminated)
	);

	step4_timer timer (
		.clk        (clk_clk),                               //   clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),   // reset.reset_n
		.address    (mm_interconnect_0_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver1_irq)               //   irq.irq
	);

	step4_mm_interconnect_0 mm_interconnect_0 (
		.CLOCK_50_clk_clk                                  (clk_clk),                                                       //                                CLOCK_50_clk.clk
		.jtag_uart_reset_reset_bridge_in_reset_reset       (rst_controller_reset_out_reset),                                //       jtag_uart_reset_reset_bridge_in_reset.reset
		.nios2_processor_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                            // nios2_processor_reset_reset_bridge_in_reset.reset
		.nios2_processor_data_master_address               (nios2_processor_data_master_address),                           //                 nios2_processor_data_master.address
		.nios2_processor_data_master_waitrequest           (nios2_processor_data_master_waitrequest),                       //                                            .waitrequest
		.nios2_processor_data_master_byteenable            (nios2_processor_data_master_byteenable),                        //                                            .byteenable
		.nios2_processor_data_master_read                  (nios2_processor_data_master_read),                              //                                            .read
		.nios2_processor_data_master_readdata              (nios2_processor_data_master_readdata),                          //                                            .readdata
		.nios2_processor_data_master_readdatavalid         (nios2_processor_data_master_readdatavalid),                     //                                            .readdatavalid
		.nios2_processor_data_master_write                 (nios2_processor_data_master_write),                             //                                            .write
		.nios2_processor_data_master_writedata             (nios2_processor_data_master_writedata),                         //                                            .writedata
		.nios2_processor_data_master_debugaccess           (nios2_processor_data_master_debugaccess),                       //                                            .debugaccess
		.nios2_processor_instruction_master_address        (nios2_processor_instruction_master_address),                    //          nios2_processor_instruction_master.address
		.nios2_processor_instruction_master_waitrequest    (nios2_processor_instruction_master_waitrequest),                //                                            .waitrequest
		.nios2_processor_instruction_master_read           (nios2_processor_instruction_master_read),                       //                                            .read
		.nios2_processor_instruction_master_readdata       (nios2_processor_instruction_master_readdata),                   //                                            .readdata
		.nios2_processor_instruction_master_readdatavalid  (nios2_processor_instruction_master_readdatavalid),              //                                            .readdatavalid
		.HEX0_s1_address                                   (mm_interconnect_0_hex0_s1_address),                             //                                     HEX0_s1.address
		.HEX0_s1_write                                     (mm_interconnect_0_hex0_s1_write),                               //                                            .write
		.HEX0_s1_readdata                                  (mm_interconnect_0_hex0_s1_readdata),                            //                                            .readdata
		.HEX0_s1_writedata                                 (mm_interconnect_0_hex0_s1_writedata),                           //                                            .writedata
		.HEX0_s1_chipselect                                (mm_interconnect_0_hex0_s1_chipselect),                          //                                            .chipselect
		.HEX1_s1_address                                   (mm_interconnect_0_hex1_s1_address),                             //                                     HEX1_s1.address
		.HEX1_s1_write                                     (mm_interconnect_0_hex1_s1_write),                               //                                            .write
		.HEX1_s1_readdata                                  (mm_interconnect_0_hex1_s1_readdata),                            //                                            .readdata
		.HEX1_s1_writedata                                 (mm_interconnect_0_hex1_s1_writedata),                           //                                            .writedata
		.HEX1_s1_chipselect                                (mm_interconnect_0_hex1_s1_chipselect),                          //                                            .chipselect
		.HEX2_s1_address                                   (mm_interconnect_0_hex2_s1_address),                             //                                     HEX2_s1.address
		.HEX2_s1_write                                     (mm_interconnect_0_hex2_s1_write),                               //                                            .write
		.HEX2_s1_readdata                                  (mm_interconnect_0_hex2_s1_readdata),                            //                                            .readdata
		.HEX2_s1_writedata                                 (mm_interconnect_0_hex2_s1_writedata),                           //                                            .writedata
		.HEX2_s1_chipselect                                (mm_interconnect_0_hex2_s1_chipselect),                          //                                            .chipselect
		.HEX3_s1_address                                   (mm_interconnect_0_hex3_s1_address),                             //                                     HEX3_s1.address
		.HEX3_s1_write                                     (mm_interconnect_0_hex3_s1_write),                               //                                            .write
		.HEX3_s1_readdata                                  (mm_interconnect_0_hex3_s1_readdata),                            //                                            .readdata
		.HEX3_s1_writedata                                 (mm_interconnect_0_hex3_s1_writedata),                           //                                            .writedata
		.HEX3_s1_chipselect                                (mm_interconnect_0_hex3_s1_chipselect),                          //                                            .chipselect
		.HEX4_s1_address                                   (mm_interconnect_0_hex4_s1_address),                             //                                     HEX4_s1.address
		.HEX4_s1_write                                     (mm_interconnect_0_hex4_s1_write),                               //                                            .write
		.HEX4_s1_readdata                                  (mm_interconnect_0_hex4_s1_readdata),                            //                                            .readdata
		.HEX4_s1_writedata                                 (mm_interconnect_0_hex4_s1_writedata),                           //                                            .writedata
		.HEX4_s1_chipselect                                (mm_interconnect_0_hex4_s1_chipselect),                          //                                            .chipselect
		.HEX5_s1_address                                   (mm_interconnect_0_hex5_s1_address),                             //                                     HEX5_s1.address
		.HEX5_s1_write                                     (mm_interconnect_0_hex5_s1_write),                               //                                            .write
		.HEX5_s1_readdata                                  (mm_interconnect_0_hex5_s1_readdata),                            //                                            .readdata
		.HEX5_s1_writedata                                 (mm_interconnect_0_hex5_s1_writedata),                           //                                            .writedata
		.HEX5_s1_chipselect                                (mm_interconnect_0_hex5_s1_chipselect),                          //                                            .chipselect
		.jtag_uart_avalon_jtag_slave_address               (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),         //                 jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write                 (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),           //                                            .write
		.jtag_uart_avalon_jtag_slave_read                  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),            //                                            .read
		.jtag_uart_avalon_jtag_slave_readdata              (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),        //                                            .readdata
		.jtag_uart_avalon_jtag_slave_writedata             (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),       //                                            .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest           (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest),     //                                            .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect            (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),      //                                            .chipselect
		.LEDR_s1_address                                   (mm_interconnect_0_ledr_s1_address),                             //                                     LEDR_s1.address
		.LEDR_s1_write                                     (mm_interconnect_0_ledr_s1_write),                               //                                            .write
		.LEDR_s1_readdata                                  (mm_interconnect_0_ledr_s1_readdata),                            //                                            .readdata
		.LEDR_s1_writedata                                 (mm_interconnect_0_ledr_s1_writedata),                           //                                            .writedata
		.LEDR_s1_chipselect                                (mm_interconnect_0_ledr_s1_chipselect),                          //                                            .chipselect
		.nios2_processor_debug_mem_slave_address           (mm_interconnect_0_nios2_processor_debug_mem_slave_address),     //             nios2_processor_debug_mem_slave.address
		.nios2_processor_debug_mem_slave_write             (mm_interconnect_0_nios2_processor_debug_mem_slave_write),       //                                            .write
		.nios2_processor_debug_mem_slave_read              (mm_interconnect_0_nios2_processor_debug_mem_slave_read),        //                                            .read
		.nios2_processor_debug_mem_slave_readdata          (mm_interconnect_0_nios2_processor_debug_mem_slave_readdata),    //                                            .readdata
		.nios2_processor_debug_mem_slave_writedata         (mm_interconnect_0_nios2_processor_debug_mem_slave_writedata),   //                                            .writedata
		.nios2_processor_debug_mem_slave_byteenable        (mm_interconnect_0_nios2_processor_debug_mem_slave_byteenable),  //                                            .byteenable
		.nios2_processor_debug_mem_slave_waitrequest       (mm_interconnect_0_nios2_processor_debug_mem_slave_waitrequest), //                                            .waitrequest
		.nios2_processor_debug_mem_slave_debugaccess       (mm_interconnect_0_nios2_processor_debug_mem_slave_debugaccess), //                                            .debugaccess
		.onchip_memory_s1_address                          (mm_interconnect_0_onchip_memory_s1_address),                    //                            onchip_memory_s1.address
		.onchip_memory_s1_write                            (mm_interconnect_0_onchip_memory_s1_write),                      //                                            .write
		.onchip_memory_s1_readdata                         (mm_interconnect_0_onchip_memory_s1_readdata),                   //                                            .readdata
		.onchip_memory_s1_writedata                        (mm_interconnect_0_onchip_memory_s1_writedata),                  //                                            .writedata
		.onchip_memory_s1_byteenable                       (mm_interconnect_0_onchip_memory_s1_byteenable),                 //                                            .byteenable
		.onchip_memory_s1_chipselect                       (mm_interconnect_0_onchip_memory_s1_chipselect),                 //                                            .chipselect
		.onchip_memory_s1_clken                            (mm_interconnect_0_onchip_memory_s1_clken),                      //                                            .clken
		.SW_s1_address                                     (mm_interconnect_0_sw_s1_address),                               //                                       SW_s1.address
		.SW_s1_readdata                                    (mm_interconnect_0_sw_s1_readdata),                              //                                            .readdata
		.timer_s1_address                                  (mm_interconnect_0_timer_s1_address),                            //                                    timer_s1.address
		.timer_s1_write                                    (mm_interconnect_0_timer_s1_write),                              //                                            .write
		.timer_s1_readdata                                 (mm_interconnect_0_timer_s1_readdata),                           //                                            .readdata
		.timer_s1_writedata                                (mm_interconnect_0_timer_s1_writedata),                          //                                            .writedata
		.timer_s1_chipselect                               (mm_interconnect_0_timer_s1_chipselect)                          //                                            .chipselect
	);

	step4_irq_mapper irq_mapper (
		.clk           (clk_clk),                            //       clk.clk
		.reset         (rst_controller_001_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.sender_irq    (nios2_processor_irq_irq)             //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                            // reset_in0.reset
		.reset_in1      (nios2_processor_debug_reset_request_reset), // reset_in1.reset
		.clk            (clk_clk),                                   //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),        // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req),    //          .reset_req
		.reset_req_in0  (1'b0),                                      // (terminated)
		.reset_req_in1  (1'b0),                                      // (terminated)
		.reset_in2      (1'b0),                                      // (terminated)
		.reset_req_in2  (1'b0),                                      // (terminated)
		.reset_in3      (1'b0),                                      // (terminated)
		.reset_req_in3  (1'b0),                                      // (terminated)
		.reset_in4      (1'b0),                                      // (terminated)
		.reset_req_in4  (1'b0),                                      // (terminated)
		.reset_in5      (1'b0),                                      // (terminated)
		.reset_req_in5  (1'b0),                                      // (terminated)
		.reset_in6      (1'b0),                                      // (terminated)
		.reset_req_in6  (1'b0),                                      // (terminated)
		.reset_in7      (1'b0),                                      // (terminated)
		.reset_req_in7  (1'b0),                                      // (terminated)
		.reset_in8      (1'b0),                                      // (terminated)
		.reset_req_in8  (1'b0),                                      // (terminated)
		.reset_in9      (1'b0),                                      // (terminated)
		.reset_req_in9  (1'b0),                                      // (terminated)
		.reset_in10     (1'b0),                                      // (terminated)
		.reset_req_in10 (1'b0),                                      // (terminated)
		.reset_in11     (1'b0),                                      // (terminated)
		.reset_req_in11 (1'b0),                                      // (terminated)
		.reset_in12     (1'b0),                                      // (terminated)
		.reset_req_in12 (1'b0),                                      // (terminated)
		.reset_in13     (1'b0),                                      // (terminated)
		.reset_req_in13 (1'b0),                                      // (terminated)
		.reset_in14     (1'b0),                                      // (terminated)
		.reset_req_in14 (1'b0),                                      // (terminated)
		.reset_in15     (1'b0),                                      // (terminated)
		.reset_req_in15 (1'b0)                                       // (terminated)
	);

endmodule
