
module step5 (
	clk_clk,
	ledr_export,
	prime_number_readdata,
	reset_reset_n);	

	input		clk_clk;
	output	[9:0]	ledr_export;
	output	[31:0]	prime_number_readdata;
	input		reset_reset_n;
endmodule
